// -----------------------------------------------------------------------------
// Copyright (c) 2014-2019 All rights reserved
// -----------------------------------------------------------------------------
// Author : Javen   penguinleo@163.com
// File   : ShiftRegister_Rx.v
// Create : 2019-11-26 16:53:42
// Revise : 2019-11-26 16:53:42
// Editor : sublime text3, tab size (4)
// Comment: this module is designed to receive the serial data and save it as byte data
//          the acquisition frequent is 16 times of baudrate, and the acquisition signal 
//          was generated by the the baudrate module.
//          The acquisition result is the 7th acquisition point, consider a better acqui-
//          -sition method, simple and reliable
//          2019-12-18   
//              The shift register is controlling the state machine during bit time. The 
//          width counter register is acting as a synchronous divider of the acquisition 
//          signal. The counter should be synchronoused with the Rx signal and count the 
//          acquisition signal. The baudrate detection and bit error detection are reali-
//          -zed in this module. And this module generate the trigger signal for the Par-
//          -ityGenerator module, FSM_Rx module, ByteAnalyse module.
//              In this module all register should be freshed synchronously with the ac-
//          -quisiiotn signal. But the falling edge of the Rx is not synchronous with the 
//          acquisition signal, the reset of the state machine and the bit width control
//          is controlled by this signal. 
//          Up module:
//              RxCore.v
//          Sub module:
//              ----
// Input Signal List:
//      1   |   clk             :   clock signal
//      2   |   rst             :   reset signal
//      3   |   AcqSig_i        :   The acquisition signal, this signal is generated by the BaudrateModule
//                                  which is designed 16 times of baudrate signal
//      4   |   Rx_i            :   The received signal which is asynchronous signal and should be synchronoused
//      5   |   State_i         :   Single hot code state code design
//      6   |   ParityResult_i  :   The parity calculate result, the parity generate module would give out the p-
//                                  -arity result at 1 clock after the 8th data bit is acquisited by the shift 
//                                  register module.
// Output Signal List:
//      1   |   BitWidthCnt_o   :   The bit width counter register, which is counting the acquisition signal to 
//                                  determine the acquisition point, the register fresh time point, and check the 
//                                  baudrate precision of the receiving signal.
//                                  The counter would start at 1 and gain to 15 then 0, next start another bit r-
//                                  -eceiving.
//      2   |   Byte_o          :   The reveiving byte from the rx wire, the byte including the start bit, data bits,
//                                  parity bits(if enabled), stop bit.
//      3   |   Bit_Synch_o     :   The synchronous signal for bit. During the last acquision signal period, this 
//                                  signal would keep high, which means next period is a new bit.
//      4   |   Rx_Synch_o      :   It is an important sychronous signal, which sychronous the RxCore with the input 
//                                  rx signal.
// Note:    2019-12-02
//              1   |   Prob1   |   The bit_width_cnt_r is better to be reinforced by tri-mode redundancy design;
//              2   |   Prob2   |   The byte_r is better to be reinforced by tri-mode redundancy design;
//          2019-12-03
//              1   |   Prob3   |   The Bit_Synch_o signal is trigger signal for the FSM, it is an important signal;
//          2019-12-04
//              1   |   Prob4   |   The FIFO write opperation is better to be inserted into the shiftresigter module;
//          2019-12-14
//              1   |   Ans_4   |   Consider agian the Prob4 should be applied in other module! 
//                                  The parity result bits was added into the byte_r, after the parity bits
//          2019-12-17
//              1   |   Prob5   |   The shift register maybe wrong, the shift register would fresh at each clock, while
//                                  the judgement would last a long time, many many clocks, it is a serious problem, the 
//                                  shift register byte_r would change many times during the judgement is available.
// -----------------------------------------------------------------------------
module ShiftRegister_Rx(
    // System signal definition
        input           clk,
        input           rst,
    // the interface with the BaudrateModule
        input           AcqSig_i,
    // the interface of the RX core
        input           Rx_i,
    // the interface with the FSM_Rx module
        input   [4:0]   State_i,
        output  [3:0]   BitWidthCnt_o,   // the index of the bit in the byte
    // the interface with the parity generator module
        input           ParityResult_i,
    // the output of the module
        output  [11:0]  Byte_o,     // the output of the shift register, including the data bits and the parity bit
    // the sychronization signal
        output          Bit_Synch_o, // a bit has been received,the bit width counter has finished
        output          Rx_Synch_o, // at the falling edge of the RX when the state machine is idle
        output          p_ParityCalTrigger_o  // the signal trigger the parity generate module
    );
    // register definition
        reg [2:0]   shift_acq_r;        // the acquisition signal delay register
        reg [2:0]   shift_reg_r;        // synchronousing the asynchronous signal 
        reg [15:0]  serial_reg_r;
        reg [3:0]   bit_width_cnt_r;   // this register was applied to measure the width of the rx signal 
        reg [11:0]  byte_r;             // this register is working like a shift register
        reg         parity_error_r;     // the parity fail
    // wire definition 
        wire        falling_edge_rx_w;  // the falling edge of the rx port
        wire        acqsig_dly_1clk_w;  // the AcqSig_i delay 1 clock output
        wire        acqsig_dly_2clk_w;  // the AcqSig_i delay 2 clock output
        wire        acqsig_dly_3clk_w;  // the AcqSig_i delay 3 clock output
    // parameter definition
        // Receiving state machine definition  
            parameter   IDLE        = 5'b0_0001;   
            parameter   STARTBIT    = 5'b0_0010;
            parameter   DATABITS    = 5'b0_0100;
            parameter   PARITYBIT   = 5'b0_1000;
            parameter   STOPBIT     = 5'b1_0000;
        // the acquisition point definition
            parameter   ACQSITION_POINT = 4'd7;
            // parameter   PARITY_POINT    = ACQSITION_POINT + 1'b1;
        // error definition
            parameter   WRONG       = 1'b1;
            parameter   RIGHT       = 1'b0;  
    // wire assign 
        assign falling_edge_rx_w    = shift_reg_r[2] & !shift_reg_r[1]; // falling edge of the rx
        assign acqsig_dly_1clk_w    = shift_acq_r[0];
        assign acqsig_dly_2clk_w    = shift_acq_r[1];
        assign acqsig_dly_3clk_w    = shift_acq_r[2];
        assign Rx_Synch_o           = falling_edge_rx_w & (State_i == IDLE);
        assign Bit_Synch_o          = ~(bit_width_cnt_r[0] | bit_width_cnt_r[1] | bit_width_cnt_r[2] | bit_width_cnt_r[3]);
        assign Byte_o               = byte_r;
        assign BitWidthCnt_o        = bit_width_cnt_r;
        assign p_ParityCalTrigger_o = (State_i == DATABITS) & (bit_width_cnt_r == ACQSITION_POINT) & (acqsig_dly_2clk_w == 1'b1); // this design each data bit freshing the parity result
    // Shift register for AcqSig_i delay
        always @(posedge clk or negedge rst) begin
            if (!rst) begin
                shift_acq_r <= 3'b000;
            end
            else begin
                shift_acq_r <= {shift_acq_r[1:0],AcqSig_i};
            end
        end
    // Shift register operation definition
        always @(posedge clk or negedge rst) begin
            if (!rst) begin
                shift_reg_r <= 3'b000;            
            end
            else if (AcqSig_i == 1'b1) begin
                shift_reg_r <= {shift_reg_r[1:0],Rx_i};
            end
            else begin
                shift_reg_r <= shift_reg_r;
            end
        end
    // serial data register operation  *the acquisition point* 
        always @(posedge clk or negedge rst) begin
            if (!rst) begin
                serial_reg_r <= 16'd0;                
            end
            else if (AcqSig_i == 1'b1) begin
                serial_reg_r <= {serial_reg_r[14:0],shift_reg_r[2]};
            end
            else begin
                serial_reg_r <= serial_reg_r;
            end
        end
    // bit width counter,Once the system was synchronized the counter is started until the end of the byte
        always @(posedge clk or negedge rst) begin   
            if (!rst) begin
                bit_width_cnt_r <= 4'd0;                
            end
            else if ((State_i == IDLE) && (falling_edge_rx_w == 1'd0) && (AcqSig_i == 1'b1)) begin
                bit_width_cnt_r <= 4'd0;
            end
            else if (Rx_Synch_o == 1'b1 && (AcqSig_i == 1'b1)) begin // equivalent to (State_i == IDLE) && (falling_edge_rx_w == 1'd1)
                bit_width_cnt_r <= 4'd1;
            end
            else if ((State_i != IDLE) && (AcqSig_i == 1'b1)) begin
                bit_width_cnt_r <= bit_width_cnt_r + 1'b1;
            end
            else begin
                bit_width_cnt_r <= bit_width_cnt_r;
            end
        end
    // byte register refresh
        always @(posedge clk or negedge rst) begin
            if (!rst) begin
                byte_r <= 12'b0000_0000_0000;                
            end
            else if ((State_i == IDLE)) begin
                byte_r <= 12'b0000_0000_0000;
            end
            else if ((State_i == STARTBIT) && (bit_width_cnt_r == ACQSITION_POINT) && (acqsig_dly_1clk_w == 1'b1)) begin   // the start bit
                byte_r <= {byte_r[10:0],shift_reg_r[2]};
            end
            else if ((State_i == DATABITS) && (bit_width_cnt_r == ACQSITION_POINT) && (acqsig_dly_1clk_w == 1'b1)) begin   // the data bits
                byte_r <= {byte_r[10:0],shift_reg_r[2]};
            end
            else if ((State_i == PARITYBIT) && (bit_width_cnt_r == ACQSITION_POINT) && (acqsig_dly_3clk_w == 1'b1)) begin  // the parity bit if the FSM move to this state
                byte_r <= {byte_r[9:0],shift_reg_r[2],ParityResult_i};  // at this point the parity calculated by this module and received parity bit are all ready
            end
            else if ((State_i == STOPBIT) && (bit_width_cnt_r == ACQSITION_POINT) && (acqsig_dly_1clk_w == 1'b1)) begin    // the stop bit
                byte_r <= {byte_r[10:0],shift_reg_r[2]};
            end
            else begin
                byte_r <= byte_r;
            end
        end
endmodule
